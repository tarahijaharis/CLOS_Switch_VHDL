LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY switch_2x2 IS
PORT	 (
	X: IN STD_LOGIC_VECTOR(7 downto 0);
	Y: IN STD_LOGIC_VECTOR(7 downto 0);
	S: IN STD_LOGIC;
	U: OUT STD_LOGIC_VECTOR(7 downto 0);
	V: OUT STD_LOGIC_VECTOR(7 downto 0)
);
END switch_2x2;

ARCHITECTURE arch_switch_2x2 OF switch_2x2 IS 
BEGIN
	U <= X WHEN S = '0' ELSE Y;
	V <= Y WHEN S = '0' ELSE X;
END ARCHITECTURE;